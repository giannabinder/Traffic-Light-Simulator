library ieee;
use ieee.std_logic_1164.all;


entity synchronizer is port (

			clk					: in std_logic;
			reset					: in std_logic;
			din					: in std_logic;
			dout					: out std_logic
  );
 end synchronizer;
 
 
architecture circuit of synchronizer is

	--component DFF_circuit is port (

			--clk					: in std_logic;
			--reset					: in std_logic;
			--d					   : in std_logic;
			--q   					: out std_logic
	  --);
	 --end component;

	Signal sreg				: std_logic_vector(1 downto 0);

BEGIN

	process(clk, reset)
	begin
		if (reset = '1') then
			sreg <= "00";
		
		elsif (rising_edge(clk)) then
			sreg(1) <= sreg(0);
			sreg(0) <= din;
		end if;
		
		dout <= sreg(1);
		
	end process;

	--inst1: DFF_circuit port map(clk, reset, din, sreg);
	--inst2: DFF_circuit port map(clk, reset, sreg, dout);
	
	

end circuit;